master \$1 $1 ( , [$1] <> slave )

