control $1 \$1 (,[$1] <> worker)
