#!/helios/bin/cdl
master \$1 \$2 [$1] ||| worker
