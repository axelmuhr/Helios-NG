#! cdl

control $1 <> ( | [i < $1] (worker %i $1))

