#! cdl

control <> ( | [$1] worker)

