#! cdl

component ccontrol { code ../pi_ring/control; }
component cworker  { code ../pi_ring/worker; }
component fworker  { code ../pi_fort/worker; }
component pworker  { code ../pi_pasc/worker; }

ccontrol <> ( (| [$1] cworker) | (| [$2] fworker) | (| [$3] pworker) )


